// perf.v - Performance Monitors for ACCEL-v1
// MAC utilization, reuse metrics, roofline
// Implements counters and roofline metrics for reuse and efficiency

// TODO: Implement performance monitoring hardware
module perf_monitor (
    // TODO: Add interface
);

endmodule