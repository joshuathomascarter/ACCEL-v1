// dma_lite.v - DMA Engine for ACCEL-v1
// AXI-Stream DMA-lite for BRAM transfers
// Implements burst DMA controller for high-bandwidth transfer

// TODO: Implement DMA lite engine
module dma_lite (
    // TODO: Add AXI-Stream interface
);

endmodule